module bridge(input clk, INF.bridge_inf inf);



endmodule