
module OS(input clk, INF.OS_inf inf);
import usertype::*;
//===========================================================================
// local parameter
//===========================================================================

//===========================================================================
// FSM
//===========================================================================

//===========================================================================
// design
//===========================================================================





//===========================================================================
// output
//===========================================================================



endmodule